
module inv
	(input x, 
	 output y);
	
	assign y = ~x;

endmodule 